//-- Megaherzios  MHz
`define F_4MHz 3
`define F_1MHz 12
    
//-- Hertzios (Hz)
`define F_2Hz   6_000_000
`define F_1Hz   12_000_000
